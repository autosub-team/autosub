
ARCHITECTURE behavior OF timingDemo IS

BEGIN
  p1 : PROCESS() --add sesitivity list for the signal connecting to port E
	--remeber to creat a variable here
   BEGIN



   END PROCESS;


 p2: PROCESS() --add sesitivity list for the signals connecting to port O and port P
  BEGIN


  END PROCESS;
--transmit the signal to the port
	N<=;
	O<=;
	P<=;
	E<=;
END behavior;

library IEEE;
use IEEE.std_logic_1164.all;

architecture behavior of truth_table is

begin

end behavior;

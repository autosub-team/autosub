library IEEE;
use IEEE.std_logic_1164.all;

ENTITY timingDemo IS 
	PORT( N,O,P,E : inout integer);
END timingDemo;  

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity {{ task_name }}_tb is
end {{ task_name }}_tb;

architecture behavior of {{ task_name }}_tb is
    --put your code here
end behavior;

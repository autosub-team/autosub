library ieee;
use ieee.std_logic_1164.all;


--##########################
--######## AND GATES #######
--##########################    
    entity AND2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity AND2;

library ieee;
use ieee.std_logic_1164.all;

    entity AND3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity AND3;

library ieee;
use ieee.std_logic_1164.all;

    entity AND4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity AND4;

--##########################
--######## NAND GATES ######
--##########################    

library ieee;
use ieee.std_logic_1164.all;

    entity NAND2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity NAND2;

library ieee;
use ieee.std_logic_1164.all;

    entity NAND3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity NAND3;

library ieee;
use ieee.std_logic_1164.all;

    entity NAND4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity NAND4;

--##########################
--######## OR GATES ########
--##########################    
library ieee;
use ieee.std_logic_1164.all;

    entity OR2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity OR2;

library ieee;
use ieee.std_logic_1164.all;

    entity OR3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity OR3;

library ieee;
use ieee.std_logic_1164.all;

    entity OR4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity OR4;

--##########################
--######## NOR GATES #######
--########################## 
library ieee;
use ieee.std_logic_1164.all;   
    entity NOR2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity NOR2;

library ieee;
use ieee.std_logic_1164.all;

    entity NOR3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity NOR3;

library ieee;
use ieee.std_logic_1164.all;

    entity NOR4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity NOR4;

--##########################
--######## XOR GATES #######
--##########################  
library ieee;
use ieee.std_logic_1164.all;
  
    entity XOR2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity XOR2;

library ieee;
use ieee.std_logic_1164.all;

    entity XOR3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity XOR3;

library ieee;
use ieee.std_logic_1164.all;

    entity XOR4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity XOR4;

--##########################
--######## XNOR GATES ######
--##########################    
library ieee;
use ieee.std_logic_1164.all;

    entity XNOR2 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            O   :out std_logic
        );
    end entity XNOR2;

library ieee;
use ieee.std_logic_1164.all;

    entity XNOR3 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            O   :out std_logic
        );
    end entity XNOR3;

library ieee;
use ieee.std_logic_1164.all;

    entity XNOR4 is
        port
        (
            I1  :in  std_logic;
            I2  :in  std_logic;
            I3  :in  std_logic;
            I4  :in  std_logic;
            O   :out std_logic
        );
    end entity XNOR4;

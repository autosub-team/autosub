library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

architecture behavioral of SC_CU_beh is	

begin

end behavioral;

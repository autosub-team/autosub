library IEEE;
use IEEE.std_logic_1164.all;

entity truth_table is
    port(   A,B,C,D : in    std_logic;
            O       : out   std_logic);
end truth_table;               

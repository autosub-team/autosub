package fsm_pkg is 
   type fsm_state is 
   (
      START,
      S0,
      S1,
      S2,
      S3      
   );
end package fsm_pkg;

library IEEE;
use IEEE.std_logic_1164.all;
use work.fsm_pkg.all;

architecture behavior of fsm is

begin

end behavior;

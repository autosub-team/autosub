library IEEE;
use IEEE.std_logic_1164.all;

architecture behavior of arithmetic is

begin

end behavior;

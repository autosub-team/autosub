library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

architecture behavioral of register_file_beh is	

begin

end behavioral;

library IEEE;
use IEEE.std_logic_1164.all;

entity pwm is
    port(   CLK    : in    std_logic;
            O      : out   std_logic);
end pwm;     

library IEEE;
use IEEE.std_logic_1164.all;

architecture behavior of ROM is

begin

end behavior;
